`define TEST
